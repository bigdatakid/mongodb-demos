    "reviewDate": {
      "$date": "2016-03-18T00:00:00.000Z"
    },
    "reviewTitle": "Thin walls and crowded parking lot.",
    "reviewText": "Hotel was ok but very thin walls - could hear conversation of room next door and people kept us up all night. The parking lot was very crowded and not well lit far away from hotel where we had to park-- was kinda scary to walk thru at night. Room was clean and spacey just too thin walls",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 3
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-02-18T00:00:00.000Z"
    },
    "reviewTitle": "Thin walls and crowded parking lot.",
    "reviewText": "Averagely nice..",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 4
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-07-22T00:00:00.000Z"
    },
    "reviewTitle": "Concert Night Stay",
    "reviewText": "Enjoyed our stay despite the fact the front desk clerk could not find our reservation when we first got there. But once I called Hotels.Com they called the hotel and resolved the problem immediately!",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 5
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2015-10-12T00:00:00.000Z"
    },
    "reviewTitle": "an expensive Austin hotel",
    "reviewText": "disappointing (370 for 2 nights - breakfast not included, shower handle broken, lavatory wouldn't drain properly (called housekeeping, but the guy didn't fix either)), could not control ac fan speed (either it was off or going full blast).",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 2
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-02-26T00:00:00.000Z"
    },
    "reviewTitle": "an expensive Austin hotel",
    "reviewText": "They said thr will be 2 complimentry water bottel en the room and thr was nothing that sucks",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 3
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-06-17T00:00:00.000Z"
    },
    "reviewTitle": "Last minute stay",
    "reviewText": "My visit was very last minute. I checked in at 10:30pm and checked out at 11:30am the following day. It was clean and comfortable. There was a side pantry downstairs for late night snacking but few healthy options. There is an all you can eat breakfast in the morning for close to 11.",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 4
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-10-28T00:00:00.000Z"
    },
    "reviewTitle": "Clean hotel and helpful staff!",
    "reviewText": "Hotel staff were amazing!! They went above and beyond to help us find great places to eat and things to do!! So nice!! Thanks so much!!",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 5
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2015-08-10T00:00:00.000Z"
    },
    "reviewTitle": "Clean hotel and helpful staff!",
    "reviewText": "Awesome hotel, very clean .... . .. ... .. ... ...............,,,,,,,,,,,,,,,,,",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 5
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-10-01T00:00:00.000Z"
    },
    "reviewTitle": "Nice over all, good place and a good value",
    "reviewText": "Good",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 4
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-01-14T00:00:00.000Z"
    },
    "reviewTitle": "Nice over all, good place and a good value",
    "reviewText": "Hotel in renovations. It isn't even old. But the rooms smelled like strong sweat and mildew. Had to move rooms from 1st floor to 2nd. Still smelled. Assuming it had to do with flooring or renovations. Otherwise it was great. Nice hotel, good breakfast and decor inside and windows. Bathrooms could have better lighting and nicer shower.",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 3
  }, {
    "reviewId": "",
