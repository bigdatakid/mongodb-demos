    "reviewText": "Nice place and shopping, eating near hotel. Everything OK. Easy to go everywhere.",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 5
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-06-30T00:00:00.000Z"
    },
    "reviewTitle": "Good for one night",
    "reviewText": "The hotel is right next to I-10 so was very convenient for one night on a road trip. The room is modern and comfortable but the breakfast was one of the poorest offerings for similarly priced hotels.",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 3
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-07-07T00:00:00.000Z"
    },
    "reviewTitle": "Good hotel, good service. Thank you.",
    "reviewText": "N/A",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 5
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-06-29T00:00:00.000Z"
    },
    "reviewTitle": "Good hotel, good service. Thank you.",
    "reviewText": "Dirty room with cokroch in bed , hair all over the place ,don't stay here",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 1
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2015-09-15T00:00:00.000Z"
    },
    "reviewTitle": "New management...great experience!!!",
    "reviewText": "I stayed here for 2 nights and paid only 92 although it still would have been worth it to pay more. I didn't expect for this place to be so clean and updated since it was cheap but I was pleasantly surprised. Everything at this hotel was spotless and the room was very nice and accommodating. I was able to do a load of laundry for 2 and it was nice to have a continental breakfast and coffee to start my day. Along with their high standards of taking care of their rooms and property in general, they have a very friendly and positive group of employees. The staff was very friendly and helpful with every question I had and constantly smiling and greeting everyone that came through their door. The manager of the hotel even offered to give me a ride to the Greyhound bus station since I checked out at 12 and didn't leave until 5pm. This place went above and beyond to make me feel comfortable and welcome. Everytime I come to El Paso I will definitely be staying here and I would recommend it to everyone traveling through here.",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 5
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2015-09-05T00:00:00.000Z"
    },
    "reviewTitle": "Great stay at a great price!",
    "reviewText": "It was great for the price I paid",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 4
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-07-18T00:00:00.000Z"
    },
    "reviewTitle": "Ok",
    "reviewText": "It was ok",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 3
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2015-09-18T00:00:00.000Z"
    },
    "reviewTitle": "Great overall experience.",
    "reviewText": "Great location at a great price. Need more pillows!!",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 5
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-06-08T00:00:00.000Z"
    },
    "reviewTitle": "Good",
    "reviewText": "Great!",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 4
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-07-31T00:00:00.000Z"
    },
    "reviewTitle": "Ok hotel",
    "reviewText": "The hotel price was good but the room was not very clean and it smell bad",
    "reviewerCity": "",
    "reviewerState": "",
    "reviewRating": 3
  }, {
    "reviewId": "",
    "reviewDate": {
      "$date": "2016-05-31T00:00:00.000Z"
    },
    "reviewTitle": "Ok hotel",
